`timescale 1ps / 1ps
module SobelFilter_Div_31Ux3U_8U_4(
          in2,
          in1,
          out1,
          clk,
          stall
);
   input [30:0] in2;
   input [2:0] in1;
   output [7:0] out1;
   input clk;
   input stall;
wire sub_145_2_n_1, sub_145_2_n_2, sub_145_2_n_3, sub_164_2_n_0, sub_164_2_n_1,
     sub_164_2_n_2, sub_164_2_n_4, sub_183_2_n_0, sub_183_2_n_1, sub_183_2_n_2,
     sub_183_2_n_3, sub_183_2_n_5, sub_183_2_n_7, sub_202_2_n_0, sub_202_2_n_1,
     sub_202_2_n_2, sub_202_2_n_3, sub_202_2_n_5, sub_202_2_n_7, sub_221_2_n_0,
     sub_221_2_n_1, sub_221_2_n_2, sub_221_2_n_3, sub_221_2_n_5, sub_221_2_n_7,
     sub_240_2_n_0, sub_240_2_n_1, sub_240_2_n_2, sub_240_2_n_3, sub_240_2_n_5,
     sub_240_2_n_7, sub_259_2_n_0, sub_259_2_n_1, sub_259_2_n_2, sub_259_2_n_3,
     sub_259_2_n_5, sub_259_2_n_7, sub_278_2_n_0, sub_278_2_n_1, sub_278_2_n_2,
     sub_278_2_n_3, sub_278_2_n_5, sub_278_2_n_7, sub_297_2_n_0, sub_297_2_n_1,
     sub_297_2_n_2, sub_297_2_n_3, sub_297_2_n_5, sub_297_2_n_7, sub_316_2_n_0,
     sub_316_2_n_1, sub_316_2_n_2, sub_316_2_n_3, sub_316_2_n_5, sub_316_2_n_7,
     sub_335_2_n_0, sub_335_2_n_1, sub_335_2_n_2, sub_335_2_n_3, sub_335_2_n_5,
     sub_335_2_n_7, sub_354_2_n_0, sub_354_2_n_1, sub_354_2_n_2, sub_354_2_n_3,
     sub_354_2_n_5, sub_354_2_n_7, sub_373_2_n_0, sub_373_2_n_1, sub_373_2_n_2,
     sub_373_2_n_3, sub_373_2_n_5, sub_373_2_n_7, sub_392_2_n_0, sub_392_2_n_1,
     sub_392_2_n_2, sub_392_2_n_3, sub_392_2_n_5, sub_392_2_n_7, sub_411_2_n_0,
     sub_411_2_n_1, sub_411_2_n_2, sub_411_2_n_3, sub_411_2_n_5, sub_411_2_n_7,
     sub_430_2_n_0, sub_430_2_n_1, sub_430_2_n_2, sub_430_2_n_3, sub_430_2_n_5,
     sub_430_2_n_7, sub_449_2_n_0, sub_449_2_n_1, sub_449_2_n_2, sub_449_2_n_3,
     sub_449_2_n_5, sub_449_2_n_7, sub_468_2_n_0, sub_468_2_n_1, sub_468_2_n_2,
     sub_468_2_n_3, sub_468_2_n_5, sub_468_2_n_7, sub_487_2_n_0, sub_487_2_n_1,
     sub_487_2_n_2, sub_487_2_n_3, sub_487_2_n_5, sub_487_2_n_7, sub_506_2_n_0,
     sub_506_2_n_1, sub_506_2_n_2, sub_506_2_n_3, sub_506_2_n_5, sub_506_2_n_7,
     sub_525_2_n_0, sub_525_2_n_1, sub_525_2_n_2, sub_525_2_n_3, sub_525_2_n_5,
     sub_525_2_n_7, sub_544_2_n_0, sub_544_2_n_1, sub_544_2_n_2, sub_544_2_n_3,
     sub_544_2_n_5, sub_544_2_n_7, sub_563_2_n_0, sub_563_2_n_1, sub_563_2_n_2,
     sub_563_2_n_3, sub_563_2_n_5, sub_563_2_n_7, sub_582_2_n_0, sub_582_2_n_1,
     sub_582_2_n_2, sub_582_2_n_3, sub_582_2_n_5, sub_582_2_n_7, sub_603_2_n_0,
     sub_603_2_n_1, sub_603_2_n_2, sub_603_2_n_3, sub_603_2_n_5, sub_603_2_n_7,
     sub_624_2_n_0, sub_624_2_n_1, sub_624_2_n_2, sub_624_2_n_3, sub_624_2_n_5,
     sub_624_2_n_7, sub_645_2_n_0, sub_645_2_n_1, sub_645_2_n_2, sub_645_2_n_3,
     sub_645_2_n_5, sub_645_2_n_7, sub_666_2_n_0, sub_666_2_n_1, sub_666_2_n_2,
     sub_666_2_n_3, sub_666_2_n_5, sub_666_2_n_7, sub_687_2_n_0, sub_687_2_n_1,
     sub_687_2_n_2, sub_687_2_n_3, sub_687_2_n_5, sub_687_2_n_7, sub_708_2_n_0,
     sub_708_2_n_1, sub_708_2_n_2, sub_708_2_n_3, sub_708_2_n_5, sub_708_2_n_7,
     sub_727_2_n_1, sub_727_2_n_2, sub_727_2_n_3, sub_727_2_n_4, sub_727_2_n_5,
     sub_727_2_n_6, sub_727_2_n_7, stall, clk, n_28, n_29, n_30, n_31, n_32,
     n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40, n_41, asc001_0_0_,
     asc001_0_1_, asc001_0_2_, asc001_0_3_, asc001_0_4_, asc001_0_5_,
     asc001_0_6_, asc001_0_7_, in2_1_0_, in2_1_3_, in2_2_0_, in2_4_0_, in2_4_1_,
     in2_4_3_, in2_5_0_, in2_5_1_, in2_7_0_, in2_7_1_, in2_7_2_, in2_7_3_,
     in2_8_0_, in2_8_1_, in2_8_2_, in2_10_0_, in2_10_1_, in2_10_2_, in2_10_3_,
     in2_11_0_, in2_11_1_, in2_11_2_, in2_13_0_, in2_13_1_, in2_13_2_, in2_13_3_,
     in2_14_0_, in2_14_1_, in2_14_2_, in2_16_0_, in2_16_1_, in2_16_2_, in2_16_3_,
     in2_17_0_, in2_17_1_, in2_17_2_, in2_19_0_, in2_19_1_, in2_19_2_, in2_19_3_,
     in2_20_0_, in2_20_1_, in2_20_2_, in2_22_0_, in2_22_1_, in2_22_2_, in2_22_3_,
     in2_23_0_, in2_23_1_, in2_23_2_, in2_25_0_, in2_25_1_, in2_25_2_, in2_25_3_,
     in2_26_0_, in2_26_1_, in2_26_2_, in2_28_0_, in2_28_1_, in2_28_2_, in2_28_3_,
     in2_29_0_, in2_29_1_, in2_29_2_, in2_31_0_, in2_31_1_, in2_31_2_, in2_31_3_,
     in2_32_0_, in2_32_1_, in2_32_2_, in2_34_0_, in2_34_1_, in2_34_2_, in2_34_3_,
     in2_35_0_, in2_35_1_, in2_35_2_, in2_37_0_, in2_37_1_, in2_37_2_, in2_37_3_,
     in2_38_0_, in2_38_1_, in2_38_2_, in2_40_0_, in2_40_1_, in2_40_2_, in2_40_3_,
     in2_41_0_, in2_41_1_, in2_41_2_, in2_43_0_, in2_43_1_, in2_43_2_, in2_43_3_,
     in2_44_0_, in2_44_1_, in2_44_2_, in2_46_0_, in2_46_1_, in2_46_2_, in2_46_3_,
     in2_47_0_, in2_47_1_, in2_47_2_, in2_49_0_, in2_49_1_, in2_49_2_, in2_49_3_,
     in2_50_0_, in2_50_1_, in2_50_2_, in2_52_0_, in2_52_1_, in2_52_2_, in2_52_3_,
     in2_53_0_, in2_53_1_, in2_53_2_, in2_55_0_, in2_55_1_, in2_55_2_, in2_55_3_,
     in2_56_0_, in2_56_1_, in2_56_2_, in2_58_0_, in2_58_1_, in2_58_2_, in2_58_3_,
     in2_59_0_, in2_59_1_, in2_59_2_, in2_61_0_, in2_61_1_, in2_61_2_, in2_61_3_,
     in2_62_0_, in2_62_1_, in2_62_2_, in2_64_0_, in2_64_1_, in2_64_2_, in2_64_3_,
     in2_65_0_, in2_65_1_, in2_65_2_, in2_67_0_, in2_67_1_, in2_67_2_, in2_67_3_,
     in2_68_0_, in2_68_1_, in2_68_2_, in2_70_0_, in2_70_1_, in2_70_2_, in2_70_3_,
     in2_71_0_, in2_71_1_, in2_71_2_, in2_73_0_, in2_73_1_, in2_73_2_, in2_73_3_,
     in2_74_0_, in2_74_1_, in2_74_2_, in2_76_0_, in2_76_1_, in2_76_2_, in2_76_3_,
     in2_77_0_, in2_77_1_, in2_77_2_, in2_79_0_, in2_79_1_, in2_79_2_, in2_79_3_,
     in2_80_0_, in2_80_1_, in2_80_2_, in2_82_0_, in2_82_1_, in2_82_2_, in2_82_3_,
     in2_83_0_, in2_83_1_, in2_83_2_, in2_85_0_, in2_85_1_, in2_85_2_, in2_85_3_,
     in2_86_0_, in2_86_1_, in2_86_2_, in2_88_0_, in2_88_1_, in2_88_2_, in2_88_3_,
     in2_89_0_, in2_89_1_, in2_89_2_, in2_91_3_;
assign {out1[7]} = asc001_0_7_;
assign {out1[6]} = asc001_0_6_;
assign {out1[5]} = asc001_0_5_;
assign {out1[4]} = asc001_0_4_;
assign {out1[3]} = asc001_0_3_;
assign {out1[2]} = asc001_0_2_;
assign {out1[1]} = asc001_0_1_;
assign {out1[0]} = asc001_0_0_;
reg cadence_register_n_28;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_28 <= sub_727_2_n_5;
    end
 end
 assign n_28 = cadence_register_n_28;
reg cadence_register_n_29;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_29 <= in2_68_0_;
    end
 end
 assign n_29 = cadence_register_n_29;
reg cadence_register_n_30;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_30 <= in1[0];
    end
 end
 assign n_30 = cadence_register_n_30;
reg cadence_register_n_31;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_31 <= in2_68_1_;
    end
 end
 assign n_31 = cadence_register_n_31;
reg cadence_register_n_32;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_32 <= in2_68_2_;
    end
 end
 assign n_32 = cadence_register_n_32;
reg cadence_register_n_33;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_33 <= in2[5];
    end
 end
 assign n_33 = cadence_register_n_33;
reg cadence_register_n_34;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_34 <= in1[1];
    end
 end
 assign n_34 = cadence_register_n_34;
reg cadence_register_n_35;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_35 <= in2[6];
    end
 end
 assign n_35 = cadence_register_n_35;
reg cadence_register_n_36;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_36 <= in2[3];
    end
 end
 assign n_36 = cadence_register_n_36;
reg cadence_register_n_37;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_37 <= in2[4];
    end
 end
 assign n_37 = cadence_register_n_37;
reg cadence_register_n_38;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_38 <= in2[1];
    end
 end
 assign n_38 = cadence_register_n_38;
reg cadence_register_n_39;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_39 <= in2[2];
    end
 end
 assign n_39 = cadence_register_n_39;
reg cadence_register_n_40;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_40 <= in2[7];
    end
 end
 assign n_40 = cadence_register_n_40;
reg cadence_register_n_41;
 always @(posedge clk) begin
    begin
       if (stall == 1'B0) 
          cadence_register_n_41 <= in1[2];
    end
 end
 assign n_41 = cadence_register_n_41;
 assign asc001_0_0_ = ~in2_91_3_;
 assign in2_71_2_ = ((in2_70_2_ & ~in2_70_3_) | (n_31 & in2_70_3_));
 assign in2_71_1_ = ((in2_70_1_ & ~in2_70_3_) | (n_29 & in2_70_3_));
 assign in2_71_0_ = ((in2_70_0_ & ~in2_70_3_) | (n_40 & in2_70_3_));
 assign in2_68_2_ = ((in2_67_2_ & ~in2_67_3_) | (in2_65_1_ & in2_67_3_));
 assign in2_68_1_ = ((in2_67_1_ & ~in2_67_3_) | (in2_65_0_ & in2_67_3_));
 assign in2_68_0_ = ((in2_67_0_ & ~in2_67_3_) | ({in2[8]} & in2_67_3_));
 assign in2_74_2_ = ((in2_73_2_ & ~in2_73_3_) | (in2_71_1_ & in2_73_3_));
 assign in2_74_1_ = ((in2_73_1_ & ~in2_73_3_) | (in2_71_0_ & in2_73_3_));
 assign in2_74_0_ = ((in2_73_0_ & ~in2_73_3_) | (n_35 & in2_73_3_));
 assign in2_65_2_ = ((in2_64_2_ & ~in2_64_3_) | (in2_62_1_ & in2_64_3_));
 assign in2_65_1_ = ((in2_64_1_ & ~in2_64_3_) | (in2_62_0_ & in2_64_3_));
 assign in2_65_0_ = ((in2_64_0_ & ~in2_64_3_) | ({in2[9]} & in2_64_3_));
 assign in2_77_2_ = ((in2_76_2_ & ~in2_76_3_) | (in2_74_1_ & in2_76_3_));
 assign in2_77_1_ = ((in2_76_1_ & ~in2_76_3_) | (in2_74_0_ & in2_76_3_));
 assign in2_77_0_ = ((in2_76_0_ & ~in2_76_3_) | (n_33 & in2_76_3_));
 assign in2_62_2_ = ((in2_61_2_ & ~in2_61_3_) | (in2_59_1_ & in2_61_3_));
 assign in2_62_1_ = ((in2_61_1_ & ~in2_61_3_) | (in2_59_0_ & in2_61_3_));
 assign in2_62_0_ = ((in2_61_0_ & ~in2_61_3_) | ({in2[10]} & in2_61_3_));
 assign in2_80_2_ = ((in2_79_2_ & ~in2_79_3_) | (in2_77_1_ & in2_79_3_));
 assign in2_80_1_ = ((in2_79_1_ & ~in2_79_3_) | (in2_77_0_ & in2_79_3_));
 assign in2_80_0_ = ((in2_79_0_ & ~in2_79_3_) | (n_37 & in2_79_3_));
 assign in2_59_2_ = ((in2_58_2_ & ~in2_58_3_) | (in2_56_1_ & in2_58_3_));
 assign in2_59_1_ = ((in2_58_1_ & ~in2_58_3_) | (in2_56_0_ & in2_58_3_));
 assign in2_59_0_ = ((in2_58_0_ & ~in2_58_3_) | ({in2[11]} & in2_58_3_));
 assign in2_83_2_ = ((in2_82_2_ & ~in2_82_3_) | (in2_80_1_ & in2_82_3_));
 assign in2_83_1_ = ((in2_82_1_ & ~in2_82_3_) | (in2_80_0_ & in2_82_3_));
 assign in2_83_0_ = ((in2_82_0_ & ~in2_82_3_) | (n_36 & in2_82_3_));
 assign in2_56_2_ = ((in2_55_2_ & ~in2_55_3_) | (in2_53_1_ & in2_55_3_));
 assign in2_56_1_ = ((in2_55_1_ & ~in2_55_3_) | (in2_53_0_ & in2_55_3_));
 assign in2_56_0_ = ((in2_55_0_ & ~in2_55_3_) | ({in2[12]} & in2_55_3_));
 assign in2_86_2_ = ((in2_85_2_ & ~in2_85_3_) | (in2_83_1_ & in2_85_3_));
 assign in2_86_1_ = ((in2_85_1_ & ~in2_85_3_) | (in2_83_0_ & in2_85_3_));
 assign in2_86_0_ = ((in2_85_0_ & ~in2_85_3_) | (n_39 & in2_85_3_));
 assign in2_53_2_ = ((in2_52_2_ & ~in2_52_3_) | (in2_50_1_ & in2_52_3_));
 assign in2_53_1_ = ((in2_52_1_ & ~in2_52_3_) | (in2_50_0_ & in2_52_3_));
 assign in2_53_0_ = ((in2_52_0_ & ~in2_52_3_) | ({in2[13]} & in2_52_3_));
 assign in2_89_2_ = ((in2_88_2_ & ~in2_88_3_) | (in2_86_1_ & in2_88_3_));
 assign in2_89_1_ = ((in2_88_1_ & ~in2_88_3_) | (in2_86_0_ & in2_88_3_));
 assign in2_89_0_ = ((in2_88_0_ & ~in2_88_3_) | (n_38 & in2_88_3_));
 assign asc001_0_1_ = ~in2_88_3_;
 assign asc001_0_7_ = ~in2_70_3_;
 assign asc001_0_2_ = ~in2_85_3_;
 assign asc001_0_5_ = ~in2_76_3_;
 assign asc001_0_4_ = ~in2_79_3_;
 assign asc001_0_3_ = ~in2_82_3_;
 assign asc001_0_6_ = ~in2_73_3_;
 assign in2_50_2_ = ((in2_49_2_ & ~in2_49_3_) | (in2_47_1_ & in2_49_3_));
 assign in2_50_1_ = ((in2_49_1_ & ~in2_49_3_) | (in2_47_0_ & in2_49_3_));
 assign in2_50_0_ = ((in2_49_0_ & ~in2_49_3_) | ({in2[14]} & in2_49_3_));
 assign in2_47_2_ = ((in2_46_2_ & ~in2_46_3_) | (in2_44_1_ & in2_46_3_));
 assign in2_47_1_ = ((in2_46_1_ & ~in2_46_3_) | (in2_44_0_ & in2_46_3_));
 assign in2_47_0_ = ((in2_46_0_ & ~in2_46_3_) | ({in2[15]} & in2_46_3_));
 assign in2_44_2_ = ((in2_43_2_ & ~in2_43_3_) | (in2_41_1_ & in2_43_3_));
 assign in2_44_1_ = ((in2_43_1_ & ~in2_43_3_) | (in2_41_0_ & in2_43_3_));
 assign in2_44_0_ = ((in2_43_0_ & ~in2_43_3_) | ({in2[16]} & in2_43_3_));
 assign in2_41_2_ = ((in2_40_2_ & ~in2_40_3_) | (in2_38_1_ & in2_40_3_));
 assign in2_41_1_ = ((in2_40_1_ & ~in2_40_3_) | (in2_38_0_ & in2_40_3_));
 assign in2_41_0_ = ((in2_40_0_ & ~in2_40_3_) | ({in2[17]} & in2_40_3_));
 assign in2_38_2_ = ((in2_37_2_ & ~in2_37_3_) | (in2_35_1_ & in2_37_3_));
 assign in2_38_1_ = ((in2_37_1_ & ~in2_37_3_) | (in2_35_0_ & in2_37_3_));
 assign in2_38_0_ = ((in2_37_0_ & ~in2_37_3_) | ({in2[18]} & in2_37_3_));
 assign in2_35_2_ = ((in2_34_2_ & ~in2_34_3_) | (in2_32_1_ & in2_34_3_));
 assign in2_35_1_ = ((in2_34_1_ & ~in2_34_3_) | (in2_32_0_ & in2_34_3_));
 assign in2_35_0_ = ((in2_34_0_ & ~in2_34_3_) | ({in2[19]} & in2_34_3_));
 assign in2_32_2_ = ((in2_31_2_ & ~in2_31_3_) | (in2_29_1_ & in2_31_3_));
 assign in2_32_1_ = ((in2_31_1_ & ~in2_31_3_) | (in2_29_0_ & in2_31_3_));
 assign in2_32_0_ = ((in2_31_0_ & ~in2_31_3_) | ({in2[20]} & in2_31_3_));
 assign in2_29_2_ = ((in2_28_2_ & ~in2_28_3_) | (in2_26_1_ & in2_28_3_));
 assign in2_29_1_ = ((in2_28_1_ & ~in2_28_3_) | (in2_26_0_ & in2_28_3_));
 assign in2_29_0_ = ((in2_28_0_ & ~in2_28_3_) | ({in2[21]} & in2_28_3_));
 assign in2_26_2_ = ((in2_25_2_ & ~in2_25_3_) | (in2_23_1_ & in2_25_3_));
 assign in2_26_1_ = ((in2_25_1_ & ~in2_25_3_) | (in2_23_0_ & in2_25_3_));
 assign in2_26_0_ = ((in2_25_0_ & ~in2_25_3_) | ({in2[22]} & in2_25_3_));
 assign in2_23_2_ = ((in2_22_2_ & ~in2_22_3_) | (in2_20_1_ & in2_22_3_));
 assign in2_23_1_ = ((in2_22_1_ & ~in2_22_3_) | (in2_20_0_ & in2_22_3_));
 assign in2_23_0_ = ((in2_22_0_ & ~in2_22_3_) | ({in2[23]} & in2_22_3_));
 assign in2_20_2_ = ((in2_19_2_ & ~in2_19_3_) | (in2_17_1_ & in2_19_3_));
 assign in2_20_1_ = ((in2_19_1_ & ~in2_19_3_) | (in2_17_0_ & in2_19_3_));
 assign in2_20_0_ = ((in2_19_0_ & ~in2_19_3_) | ({in2[24]} & in2_19_3_));
 assign in2_17_2_ = ((in2_16_2_ & ~in2_16_3_) | (in2_14_1_ & in2_16_3_));
 assign in2_17_1_ = ((in2_16_1_ & ~in2_16_3_) | (in2_14_0_ & in2_16_3_));
 assign in2_17_0_ = ((in2_16_0_ & ~in2_16_3_) | ({in2[25]} & in2_16_3_));
 assign in2_14_2_ = ((in2_13_2_ & ~in2_13_3_) | (in2_11_1_ & in2_13_3_));
 assign in2_14_1_ = ((in2_13_1_ & ~in2_13_3_) | (in2_11_0_ & in2_13_3_));
 assign in2_14_0_ = ((in2_13_0_ & ~in2_13_3_) | ({in2[26]} & in2_13_3_));
 assign in2_11_2_ = ((in2_10_2_ & ~in2_10_3_) | (in2_8_1_ & in2_10_3_));
 assign in2_11_1_ = ((in2_10_1_ & ~in2_10_3_) | (in2_8_0_ & in2_10_3_));
 assign in2_11_0_ = ((in2_10_0_ & ~in2_10_3_) | ({in2[27]} & in2_10_3_));
 assign in2_8_2_ = ((in2_7_2_ & ~in2_7_3_) | (in2_5_1_ & in2_7_3_));
 assign in2_8_1_ = ((in2_7_1_ & ~in2_7_3_) | (in2_5_0_ & in2_7_3_));
 assign in2_8_0_ = ((in2_7_0_ & ~in2_7_3_) | ({in2[28]} & in2_7_3_));
 assign in2_5_1_ = ((in2_4_1_ & ~in2_4_3_) | (in2_2_0_ & in2_4_3_));
 assign in2_5_0_ = ((in2_4_0_ & ~in2_4_3_) | ({in2[29]} & in2_4_3_));
 assign in2_2_0_ = ((in2_1_0_ & ~in2_1_3_) | ({in2[30]} & in2_1_3_));
 assign in2_1_3_ = (sub_145_2_n_2 | ({in1[1]} | {in1[2]}));
 assign in2_1_0_ = ~sub_145_2_n_3;
 assign sub_145_2_n_2 = (sub_145_2_n_1 & {in1[0]});
 assign sub_145_2_n_3 = (sub_145_2_n_1 ^ {in1[0]});
 assign sub_145_2_n_1 = ~{in2[30]};
 assign in2_4_3_ = ~(sub_164_2_n_4 & ~{in1[2]});
 assign sub_164_2_n_4 = ((sub_164_2_n_2 & in2_2_0_) | ((in2_2_0_ & sub_164_2_n_1) | (sub_164_2_n_1 &
    sub_164_2_n_2)));
 assign in2_4_1_ = (in2_2_0_ ^ (sub_164_2_n_1 ^ sub_164_2_n_2));
 assign in2_4_0_ = ~(sub_164_2_n_2 & ~(sub_164_2_n_0 & {in2[29]}));
 assign sub_164_2_n_2 = ~({in1[0]} & ~{in2[29]});
 assign sub_164_2_n_1 = ~{in1[1]};
 assign sub_164_2_n_0 = ~{in1[0]};
 assign in2_7_3_ = ~sub_183_2_n_7;
 assign sub_183_2_n_7 = ((sub_183_2_n_5 & sub_183_2_n_0) | ((sub_183_2_n_0 & in2_5_1_) | (in2_5_1_ &
    sub_183_2_n_5)));
 assign in2_7_2_ = (sub_183_2_n_0 ^ (in2_5_1_ ^ sub_183_2_n_5));
 assign sub_183_2_n_5 = ((sub_183_2_n_3 & in2_5_0_) | ((in2_5_0_ & sub_183_2_n_2) | (sub_183_2_n_2 &
    sub_183_2_n_3)));
 assign in2_7_1_ = (in2_5_0_ ^ (sub_183_2_n_2 ^ sub_183_2_n_3));
 assign in2_7_0_ = ~(sub_183_2_n_3 & ~(sub_183_2_n_1 & {in2[28]}));
 assign sub_183_2_n_3 = ~({in1[0]} & ~{in2[28]});
 assign sub_183_2_n_2 = ~{in1[1]};
 assign sub_183_2_n_1 = ~{in1[0]};
 assign sub_183_2_n_0 = ~{in1[2]};
 assign in2_10_3_ = ~(sub_202_2_n_7 ^ in2_8_2_);
 assign sub_202_2_n_7 = ((sub_202_2_n_5 & sub_202_2_n_0) | ((sub_202_2_n_0 & in2_8_1_) | (in2_8_1_ &
    sub_202_2_n_5)));
 assign in2_10_2_ = (sub_202_2_n_0 ^ (in2_8_1_ ^ sub_202_2_n_5));
 assign sub_202_2_n_5 = ((sub_202_2_n_3 & in2_8_0_) | ((in2_8_0_ & sub_202_2_n_1) | (sub_202_2_n_1 &
    sub_202_2_n_3)));
 assign in2_10_1_ = (in2_8_0_ ^ (sub_202_2_n_1 ^ sub_202_2_n_3));
 assign in2_10_0_ = ~(sub_202_2_n_3 & ~(sub_202_2_n_2 & {in2[27]}));
 assign sub_202_2_n_3 = ~({in1[0]} & ~{in2[27]});
 assign sub_202_2_n_2 = ~{in1[0]};
 assign sub_202_2_n_1 = ~{in1[1]};
 assign sub_202_2_n_0 = ~{in1[2]};
 assign in2_13_3_ = ~(sub_221_2_n_7 ^ in2_11_2_);
 assign sub_221_2_n_7 = ((sub_221_2_n_5 & sub_221_2_n_0) | ((sub_221_2_n_0 & in2_11_1_) | (in2_11_1_
    & sub_221_2_n_5)));
 assign in2_13_2_ = (sub_221_2_n_0 ^ (in2_11_1_ ^ sub_221_2_n_5));
 assign sub_221_2_n_5 = ((sub_221_2_n_3 & in2_11_0_) | ((in2_11_0_ & sub_221_2_n_1) | (sub_221_2_n_1
    & sub_221_2_n_3)));
 assign in2_13_1_ = (in2_11_0_ ^ (sub_221_2_n_1 ^ sub_221_2_n_3));
 assign in2_13_0_ = ~(sub_221_2_n_3 & ~(sub_221_2_n_2 & {in2[26]}));
 assign sub_221_2_n_3 = ~({in1[0]} & ~{in2[26]});
 assign sub_221_2_n_2 = ~{in1[0]};
 assign sub_221_2_n_1 = ~{in1[1]};
 assign sub_221_2_n_0 = ~{in1[2]};
 assign in2_16_3_ = ~(sub_240_2_n_7 ^ in2_14_2_);
 assign sub_240_2_n_7 = ((sub_240_2_n_5 & sub_240_2_n_0) | ((sub_240_2_n_0 & in2_14_1_) | (in2_14_1_
    & sub_240_2_n_5)));
 assign in2_16_2_ = (sub_240_2_n_0 ^ (in2_14_1_ ^ sub_240_2_n_5));
 assign sub_240_2_n_5 = ((sub_240_2_n_3 & in2_14_0_) | ((in2_14_0_ & sub_240_2_n_1) | (sub_240_2_n_1
    & sub_240_2_n_3)));
 assign in2_16_1_ = (in2_14_0_ ^ (sub_240_2_n_1 ^ sub_240_2_n_3));
 assign in2_16_0_ = ~(sub_240_2_n_3 & ~(sub_240_2_n_2 & {in2[25]}));
 assign sub_240_2_n_3 = ~({in1[0]} & ~{in2[25]});
 assign sub_240_2_n_2 = ~{in1[0]};
 assign sub_240_2_n_1 = ~{in1[1]};
 assign sub_240_2_n_0 = ~{in1[2]};
 assign in2_19_3_ = ~(sub_259_2_n_7 ^ in2_17_2_);
 assign sub_259_2_n_7 = ((sub_259_2_n_5 & sub_259_2_n_0) | ((sub_259_2_n_0 & in2_17_1_) | (in2_17_1_
    & sub_259_2_n_5)));
 assign in2_19_2_ = (sub_259_2_n_0 ^ (in2_17_1_ ^ sub_259_2_n_5));
 assign sub_259_2_n_5 = ((sub_259_2_n_3 & in2_17_0_) | ((in2_17_0_ & sub_259_2_n_1) | (sub_259_2_n_1
    & sub_259_2_n_3)));
 assign in2_19_1_ = (in2_17_0_ ^ (sub_259_2_n_1 ^ sub_259_2_n_3));
 assign in2_19_0_ = ~(sub_259_2_n_3 & ~(sub_259_2_n_2 & {in2[24]}));
 assign sub_259_2_n_3 = ~({in1[0]} & ~{in2[24]});
 assign sub_259_2_n_2 = ~{in1[0]};
 assign sub_259_2_n_1 = ~{in1[1]};
 assign sub_259_2_n_0 = ~{in1[2]};
 assign in2_22_3_ = ~(sub_278_2_n_7 ^ in2_20_2_);
 assign sub_278_2_n_7 = ((sub_278_2_n_5 & sub_278_2_n_0) | ((sub_278_2_n_0 & in2_20_1_) | (in2_20_1_
    & sub_278_2_n_5)));
 assign in2_22_2_ = (sub_278_2_n_0 ^ (in2_20_1_ ^ sub_278_2_n_5));
 assign sub_278_2_n_5 = ((sub_278_2_n_3 & in2_20_0_) | ((in2_20_0_ & sub_278_2_n_1) | (sub_278_2_n_1
    & sub_278_2_n_3)));
 assign in2_22_1_ = (in2_20_0_ ^ (sub_278_2_n_1 ^ sub_278_2_n_3));
 assign in2_22_0_ = ~(sub_278_2_n_3 & ~(sub_278_2_n_2 & {in2[23]}));
 assign sub_278_2_n_3 = ~({in1[0]} & ~{in2[23]});
 assign sub_278_2_n_2 = ~{in1[0]};
 assign sub_278_2_n_1 = ~{in1[1]};
 assign sub_278_2_n_0 = ~{in1[2]};
 assign in2_25_3_ = ~(sub_297_2_n_7 ^ in2_23_2_);
 assign sub_297_2_n_7 = ((sub_297_2_n_5 & sub_297_2_n_0) | ((sub_297_2_n_0 & in2_23_1_) | (in2_23_1_
    & sub_297_2_n_5)));
 assign in2_25_2_ = (sub_297_2_n_0 ^ (in2_23_1_ ^ sub_297_2_n_5));
 assign sub_297_2_n_5 = ((sub_297_2_n_3 & in2_23_0_) | ((in2_23_0_ & sub_297_2_n_1) | (sub_297_2_n_1
    & sub_297_2_n_3)));
 assign in2_25_1_ = (in2_23_0_ ^ (sub_297_2_n_1 ^ sub_297_2_n_3));
 assign in2_25_0_ = ~(sub_297_2_n_3 & ~(sub_297_2_n_2 & {in2[22]}));
 assign sub_297_2_n_3 = ~({in1[0]} & ~{in2[22]});
 assign sub_297_2_n_2 = ~{in1[0]};
 assign sub_297_2_n_1 = ~{in1[1]};
 assign sub_297_2_n_0 = ~{in1[2]};
 assign in2_28_3_ = ~(sub_316_2_n_7 ^ in2_26_2_);
 assign sub_316_2_n_7 = ((sub_316_2_n_5 & sub_316_2_n_0) | ((sub_316_2_n_0 & in2_26_1_) | (in2_26_1_
    & sub_316_2_n_5)));
 assign in2_28_2_ = (sub_316_2_n_0 ^ (in2_26_1_ ^ sub_316_2_n_5));
 assign sub_316_2_n_5 = ((sub_316_2_n_3 & in2_26_0_) | ((in2_26_0_ & sub_316_2_n_1) | (sub_316_2_n_1
    & sub_316_2_n_3)));
 assign in2_28_1_ = (in2_26_0_ ^ (sub_316_2_n_1 ^ sub_316_2_n_3));
 assign in2_28_0_ = ~(sub_316_2_n_3 & ~(sub_316_2_n_2 & {in2[21]}));
 assign sub_316_2_n_3 = ~({in1[0]} & ~{in2[21]});
 assign sub_316_2_n_2 = ~{in1[0]};
 assign sub_316_2_n_1 = ~{in1[1]};
 assign sub_316_2_n_0 = ~{in1[2]};
 assign in2_31_3_ = ~(sub_335_2_n_7 ^ in2_29_2_);
 assign sub_335_2_n_7 = ((sub_335_2_n_5 & sub_335_2_n_0) | ((sub_335_2_n_0 & in2_29_1_) | (in2_29_1_
    & sub_335_2_n_5)));
 assign in2_31_2_ = (sub_335_2_n_0 ^ (in2_29_1_ ^ sub_335_2_n_5));
 assign sub_335_2_n_5 = ((sub_335_2_n_3 & in2_29_0_) | ((in2_29_0_ & sub_335_2_n_1) | (sub_335_2_n_1
    & sub_335_2_n_3)));
 assign in2_31_1_ = (in2_29_0_ ^ (sub_335_2_n_1 ^ sub_335_2_n_3));
 assign in2_31_0_ = ~(sub_335_2_n_3 & ~(sub_335_2_n_2 & {in2[20]}));
 assign sub_335_2_n_3 = ~({in1[0]} & ~{in2[20]});
 assign sub_335_2_n_2 = ~{in1[0]};
 assign sub_335_2_n_1 = ~{in1[1]};
 assign sub_335_2_n_0 = ~{in1[2]};
 assign in2_34_3_ = ~(sub_354_2_n_7 ^ in2_32_2_);
 assign sub_354_2_n_7 = ((sub_354_2_n_5 & sub_354_2_n_0) | ((sub_354_2_n_0 & in2_32_1_) | (in2_32_1_
    & sub_354_2_n_5)));
 assign in2_34_2_ = (sub_354_2_n_0 ^ (in2_32_1_ ^ sub_354_2_n_5));
 assign sub_354_2_n_5 = ((sub_354_2_n_3 & in2_32_0_) | ((in2_32_0_ & sub_354_2_n_1) | (sub_354_2_n_1
    & sub_354_2_n_3)));
 assign in2_34_1_ = (in2_32_0_ ^ (sub_354_2_n_1 ^ sub_354_2_n_3));
 assign in2_34_0_ = ~(sub_354_2_n_3 & ~(sub_354_2_n_2 & {in2[19]}));
 assign sub_354_2_n_3 = ~({in1[0]} & ~{in2[19]});
 assign sub_354_2_n_2 = ~{in1[0]};
 assign sub_354_2_n_1 = ~{in1[1]};
 assign sub_354_2_n_0 = ~{in1[2]};
 assign in2_37_3_ = ~(sub_373_2_n_7 ^ in2_35_2_);
 assign sub_373_2_n_7 = ((sub_373_2_n_5 & sub_373_2_n_0) | ((sub_373_2_n_0 & in2_35_1_) | (in2_35_1_
    & sub_373_2_n_5)));
 assign in2_37_2_ = (sub_373_2_n_0 ^ (in2_35_1_ ^ sub_373_2_n_5));
 assign sub_373_2_n_5 = ((sub_373_2_n_3 & in2_35_0_) | ((in2_35_0_ & sub_373_2_n_1) | (sub_373_2_n_1
    & sub_373_2_n_3)));
 assign in2_37_1_ = (in2_35_0_ ^ (sub_373_2_n_1 ^ sub_373_2_n_3));
 assign in2_37_0_ = ~(sub_373_2_n_3 & ~(sub_373_2_n_2 & {in2[18]}));
 assign sub_373_2_n_3 = ~({in1[0]} & ~{in2[18]});
 assign sub_373_2_n_2 = ~{in1[0]};
 assign sub_373_2_n_1 = ~{in1[1]};
 assign sub_373_2_n_0 = ~{in1[2]};
 assign in2_40_3_ = ~(sub_392_2_n_7 ^ in2_38_2_);
 assign sub_392_2_n_7 = ((sub_392_2_n_5 & sub_392_2_n_0) | ((sub_392_2_n_0 & in2_38_1_) | (in2_38_1_
    & sub_392_2_n_5)));
 assign in2_40_2_ = (sub_392_2_n_0 ^ (in2_38_1_ ^ sub_392_2_n_5));
 assign sub_392_2_n_5 = ((sub_392_2_n_3 & in2_38_0_) | ((in2_38_0_ & sub_392_2_n_1) | (sub_392_2_n_1
    & sub_392_2_n_3)));
 assign in2_40_1_ = (in2_38_0_ ^ (sub_392_2_n_1 ^ sub_392_2_n_3));
 assign in2_40_0_ = ~(sub_392_2_n_3 & ~(sub_392_2_n_2 & {in2[17]}));
 assign sub_392_2_n_3 = ~({in1[0]} & ~{in2[17]});
 assign sub_392_2_n_2 = ~{in1[0]};
 assign sub_392_2_n_1 = ~{in1[1]};
 assign sub_392_2_n_0 = ~{in1[2]};
 assign in2_43_3_ = ~(sub_411_2_n_7 ^ in2_41_2_);
 assign sub_411_2_n_7 = ((sub_411_2_n_5 & sub_411_2_n_0) | ((sub_411_2_n_0 & in2_41_1_) | (in2_41_1_
    & sub_411_2_n_5)));
 assign in2_43_2_ = (sub_411_2_n_0 ^ (in2_41_1_ ^ sub_411_2_n_5));
 assign sub_411_2_n_5 = ((sub_411_2_n_3 & in2_41_0_) | ((in2_41_0_ & sub_411_2_n_1) | (sub_411_2_n_1
    & sub_411_2_n_3)));
 assign in2_43_1_ = (in2_41_0_ ^ (sub_411_2_n_1 ^ sub_411_2_n_3));
 assign in2_43_0_ = ~(sub_411_2_n_3 & ~(sub_411_2_n_2 & {in2[16]}));
 assign sub_411_2_n_3 = ~({in1[0]} & ~{in2[16]});
 assign sub_411_2_n_2 = ~{in1[0]};
 assign sub_411_2_n_1 = ~{in1[1]};
 assign sub_411_2_n_0 = ~{in1[2]};
 assign in2_46_3_ = ~(sub_430_2_n_7 ^ in2_44_2_);
 assign sub_430_2_n_7 = ((sub_430_2_n_5 & sub_430_2_n_0) | ((sub_430_2_n_0 & in2_44_1_) | (in2_44_1_
    & sub_430_2_n_5)));
 assign in2_46_2_ = (sub_430_2_n_0 ^ (in2_44_1_ ^ sub_430_2_n_5));
 assign sub_430_2_n_5 = ((sub_430_2_n_3 & in2_44_0_) | ((in2_44_0_ & sub_430_2_n_1) | (sub_430_2_n_1
    & sub_430_2_n_3)));
 assign in2_46_1_ = (in2_44_0_ ^ (sub_430_2_n_1 ^ sub_430_2_n_3));
 assign in2_46_0_ = ~(sub_430_2_n_3 & ~(sub_430_2_n_2 & {in2[15]}));
 assign sub_430_2_n_3 = ~({in1[0]} & ~{in2[15]});
 assign sub_430_2_n_2 = ~{in1[0]};
 assign sub_430_2_n_1 = ~{in1[1]};
 assign sub_430_2_n_0 = ~{in1[2]};
 assign in2_49_3_ = ~(sub_449_2_n_7 ^ in2_47_2_);
 assign sub_449_2_n_7 = ((sub_449_2_n_5 & sub_449_2_n_0) | ((sub_449_2_n_0 & in2_47_1_) | (in2_47_1_
    & sub_449_2_n_5)));
 assign in2_49_2_ = (sub_449_2_n_0 ^ (in2_47_1_ ^ sub_449_2_n_5));
 assign sub_449_2_n_5 = ((sub_449_2_n_3 & in2_47_0_) | ((in2_47_0_ & sub_449_2_n_1) | (sub_449_2_n_1
    & sub_449_2_n_3)));
 assign in2_49_1_ = (in2_47_0_ ^ (sub_449_2_n_1 ^ sub_449_2_n_3));
 assign in2_49_0_ = ~(sub_449_2_n_3 & ~(sub_449_2_n_2 & {in2[14]}));
 assign sub_449_2_n_3 = ~({in1[0]} & ~{in2[14]});
 assign sub_449_2_n_2 = ~{in1[0]};
 assign sub_449_2_n_1 = ~{in1[1]};
 assign sub_449_2_n_0 = ~{in1[2]};
 assign in2_52_3_ = ~(sub_468_2_n_7 ^ in2_50_2_);
 assign sub_468_2_n_7 = ((sub_468_2_n_5 & sub_468_2_n_0) | ((sub_468_2_n_0 & in2_50_1_) | (in2_50_1_
    & sub_468_2_n_5)));
 assign in2_52_2_ = (sub_468_2_n_0 ^ (in2_50_1_ ^ sub_468_2_n_5));
 assign sub_468_2_n_5 = ((sub_468_2_n_3 & in2_50_0_) | ((in2_50_0_ & sub_468_2_n_1) | (sub_468_2_n_1
    & sub_468_2_n_3)));
 assign in2_52_1_ = (in2_50_0_ ^ (sub_468_2_n_1 ^ sub_468_2_n_3));
 assign in2_52_0_ = ~(sub_468_2_n_3 & ~(sub_468_2_n_2 & {in2[13]}));
 assign sub_468_2_n_3 = ~({in1[0]} & ~{in2[13]});
 assign sub_468_2_n_2 = ~{in1[0]};
 assign sub_468_2_n_1 = ~{in1[1]};
 assign sub_468_2_n_0 = ~{in1[2]};
 assign in2_55_3_ = ~(sub_487_2_n_7 ^ in2_53_2_);
 assign sub_487_2_n_7 = ((sub_487_2_n_5 & sub_487_2_n_0) | ((sub_487_2_n_0 & in2_53_1_) | (in2_53_1_
    & sub_487_2_n_5)));
 assign in2_55_2_ = (sub_487_2_n_0 ^ (in2_53_1_ ^ sub_487_2_n_5));
 assign sub_487_2_n_5 = ((sub_487_2_n_3 & in2_53_0_) | ((in2_53_0_ & sub_487_2_n_1) | (sub_487_2_n_1
    & sub_487_2_n_3)));
 assign in2_55_1_ = (in2_53_0_ ^ (sub_487_2_n_1 ^ sub_487_2_n_3));
 assign in2_55_0_ = ~(sub_487_2_n_3 & ~(sub_487_2_n_2 & {in2[12]}));
 assign sub_487_2_n_3 = ~({in1[0]} & ~{in2[12]});
 assign sub_487_2_n_2 = ~{in1[0]};
 assign sub_487_2_n_1 = ~{in1[1]};
 assign sub_487_2_n_0 = ~{in1[2]};
 assign in2_58_3_ = ~(sub_506_2_n_7 ^ in2_56_2_);
 assign sub_506_2_n_7 = ((sub_506_2_n_5 & sub_506_2_n_0) | ((sub_506_2_n_0 & in2_56_1_) | (in2_56_1_
    & sub_506_2_n_5)));
 assign in2_58_2_ = (sub_506_2_n_0 ^ (in2_56_1_ ^ sub_506_2_n_5));
 assign sub_506_2_n_5 = ((sub_506_2_n_3 & in2_56_0_) | ((in2_56_0_ & sub_506_2_n_1) | (sub_506_2_n_1
    & sub_506_2_n_3)));
 assign in2_58_1_ = (in2_56_0_ ^ (sub_506_2_n_1 ^ sub_506_2_n_3));
 assign in2_58_0_ = ~(sub_506_2_n_3 & ~(sub_506_2_n_2 & {in2[11]}));
 assign sub_506_2_n_3 = ~({in1[0]} & ~{in2[11]});
 assign sub_506_2_n_2 = ~{in1[0]};
 assign sub_506_2_n_1 = ~{in1[1]};
 assign sub_506_2_n_0 = ~{in1[2]};
 assign in2_61_3_ = ~(sub_525_2_n_7 ^ in2_59_2_);
 assign sub_525_2_n_7 = ((sub_525_2_n_5 & sub_525_2_n_0) | ((sub_525_2_n_0 & in2_59_1_) | (in2_59_1_
    & sub_525_2_n_5)));
 assign in2_61_2_ = (sub_525_2_n_0 ^ (in2_59_1_ ^ sub_525_2_n_5));
 assign sub_525_2_n_5 = ((sub_525_2_n_3 & in2_59_0_) | ((in2_59_0_ & sub_525_2_n_1) | (sub_525_2_n_1
    & sub_525_2_n_3)));
 assign in2_61_1_ = (in2_59_0_ ^ (sub_525_2_n_1 ^ sub_525_2_n_3));
 assign in2_61_0_ = ~(sub_525_2_n_3 & ~(sub_525_2_n_2 & {in2[10]}));
 assign sub_525_2_n_3 = ~({in1[0]} & ~{in2[10]});
 assign sub_525_2_n_2 = ~{in1[0]};
 assign sub_525_2_n_1 = ~{in1[1]};
 assign sub_525_2_n_0 = ~{in1[2]};
 assign in2_64_3_ = ~(sub_544_2_n_7 ^ in2_62_2_);
 assign sub_544_2_n_7 = ((sub_544_2_n_5 & sub_544_2_n_0) | ((sub_544_2_n_0 & in2_62_1_) | (in2_62_1_
    & sub_544_2_n_5)));
 assign in2_64_2_ = (sub_544_2_n_0 ^ (in2_62_1_ ^ sub_544_2_n_5));
 assign sub_544_2_n_5 = ((sub_544_2_n_3 & in2_62_0_) | ((in2_62_0_ & sub_544_2_n_1) | (sub_544_2_n_1
    & sub_544_2_n_3)));
 assign in2_64_1_ = (in2_62_0_ ^ (sub_544_2_n_1 ^ sub_544_2_n_3));
 assign in2_64_0_ = ~(sub_544_2_n_3 & ~(sub_544_2_n_2 & {in2[9]}));
 assign sub_544_2_n_3 = ~({in1[0]} & ~{in2[9]});
 assign sub_544_2_n_2 = ~{in1[0]};
 assign sub_544_2_n_1 = ~{in1[1]};
 assign sub_544_2_n_0 = ~{in1[2]};
 assign in2_67_3_ = ~(sub_563_2_n_7 ^ in2_65_2_);
 assign sub_563_2_n_7 = ((sub_563_2_n_5 & sub_563_2_n_0) | ((sub_563_2_n_0 & in2_65_1_) | (in2_65_1_
    & sub_563_2_n_5)));
 assign in2_67_2_ = (sub_563_2_n_0 ^ (in2_65_1_ ^ sub_563_2_n_5));
 assign sub_563_2_n_5 = ((sub_563_2_n_3 & in2_65_0_) | ((in2_65_0_ & sub_563_2_n_1) | (sub_563_2_n_1
    & sub_563_2_n_3)));
 assign in2_67_1_ = (in2_65_0_ ^ (sub_563_2_n_1 ^ sub_563_2_n_3));
 assign in2_67_0_ = ~(sub_563_2_n_3 & ~(sub_563_2_n_2 & {in2[8]}));
 assign sub_563_2_n_3 = ~({in1[0]} & ~{in2[8]});
 assign sub_563_2_n_2 = ~{in1[0]};
 assign sub_563_2_n_1 = ~{in1[1]};
 assign sub_563_2_n_0 = ~{in1[2]};
 assign in2_70_3_ = ~(sub_582_2_n_7 ^ n_32);
 assign sub_582_2_n_7 = ((sub_582_2_n_5 & sub_582_2_n_0) | ((sub_582_2_n_0 & n_31) | (n_31 & sub_582_2_n_5)));
 assign in2_70_2_ = (sub_582_2_n_0 ^ (n_31 ^ sub_582_2_n_5));
 assign sub_582_2_n_5 = ((sub_582_2_n_3 & n_29) | ((n_29 & sub_582_2_n_1) | (sub_582_2_n_1 & sub_582_2_n_3)));
 assign in2_70_1_ = (n_29 ^ (sub_582_2_n_1 ^ sub_582_2_n_3));
 assign in2_70_0_ = ~(sub_582_2_n_3 & ~(sub_582_2_n_2 & n_40));
 assign sub_582_2_n_3 = ~(n_30 & ~n_40);
 assign sub_582_2_n_2 = ~n_30;
 assign sub_582_2_n_1 = ~n_34;
 assign sub_582_2_n_0 = ~n_41;
 assign in2_73_3_ = ~(sub_603_2_n_7 ^ in2_71_2_);
 assign sub_603_2_n_7 = ((sub_603_2_n_5 & sub_603_2_n_0) | ((sub_603_2_n_0 & in2_71_1_) | (in2_71_1_
    & sub_603_2_n_5)));
 assign in2_73_2_ = (sub_603_2_n_0 ^ (in2_71_1_ ^ sub_603_2_n_5));
 assign sub_603_2_n_5 = ((sub_603_2_n_3 & in2_71_0_) | ((in2_71_0_ & sub_603_2_n_1) | (sub_603_2_n_1
    & sub_603_2_n_3)));
 assign in2_73_1_ = (in2_71_0_ ^ (sub_603_2_n_1 ^ sub_603_2_n_3));
 assign in2_73_0_ = ~(sub_603_2_n_3 & ~(sub_603_2_n_2 & n_35));
 assign sub_603_2_n_3 = ~(n_30 & ~n_35);
 assign sub_603_2_n_2 = ~n_30;
 assign sub_603_2_n_1 = ~n_34;
 assign sub_603_2_n_0 = ~n_41;
 assign in2_76_3_ = ~(sub_624_2_n_7 ^ in2_74_2_);
 assign sub_624_2_n_7 = ((sub_624_2_n_5 & sub_624_2_n_0) | ((sub_624_2_n_0 & in2_74_1_) | (in2_74_1_
    & sub_624_2_n_5)));
 assign in2_76_2_ = (sub_624_2_n_0 ^ (in2_74_1_ ^ sub_624_2_n_5));
 assign sub_624_2_n_5 = ((sub_624_2_n_3 & in2_74_0_) | ((in2_74_0_ & sub_624_2_n_1) | (sub_624_2_n_1
    & sub_624_2_n_3)));
 assign in2_76_1_ = (in2_74_0_ ^ (sub_624_2_n_1 ^ sub_624_2_n_3));
 assign in2_76_0_ = ~(sub_624_2_n_3 & ~(sub_624_2_n_2 & n_33));
 assign sub_624_2_n_3 = ~(n_30 & ~n_33);
 assign sub_624_2_n_2 = ~n_30;
 assign sub_624_2_n_1 = ~n_34;
 assign sub_624_2_n_0 = ~n_41;
 assign in2_79_3_ = ~(sub_645_2_n_7 ^ in2_77_2_);
 assign sub_645_2_n_7 = ((sub_645_2_n_5 & sub_645_2_n_0) | ((sub_645_2_n_0 & in2_77_1_) | (in2_77_1_
    & sub_645_2_n_5)));
 assign in2_79_2_ = (sub_645_2_n_0 ^ (in2_77_1_ ^ sub_645_2_n_5));
 assign sub_645_2_n_5 = ((sub_645_2_n_3 & in2_77_0_) | ((in2_77_0_ & sub_645_2_n_1) | (sub_645_2_n_1
    & sub_645_2_n_3)));
 assign in2_79_1_ = (in2_77_0_ ^ (sub_645_2_n_1 ^ sub_645_2_n_3));
 assign in2_79_0_ = ~(sub_645_2_n_3 & ~(sub_645_2_n_2 & n_37));
 assign sub_645_2_n_3 = ~(n_30 & ~n_37);
 assign sub_645_2_n_2 = ~n_30;
 assign sub_645_2_n_1 = ~n_34;
 assign sub_645_2_n_0 = ~n_41;
 assign in2_82_3_ = ~(sub_666_2_n_7 ^ in2_80_2_);
 assign sub_666_2_n_7 = ((sub_666_2_n_5 & sub_666_2_n_0) | ((sub_666_2_n_0 & in2_80_1_) | (in2_80_1_
    & sub_666_2_n_5)));
 assign in2_82_2_ = (sub_666_2_n_0 ^ (in2_80_1_ ^ sub_666_2_n_5));
 assign sub_666_2_n_5 = ((sub_666_2_n_3 & in2_80_0_) | ((in2_80_0_ & sub_666_2_n_1) | (sub_666_2_n_1
    & sub_666_2_n_3)));
 assign in2_82_1_ = (in2_80_0_ ^ (sub_666_2_n_1 ^ sub_666_2_n_3));
 assign in2_82_0_ = ~(sub_666_2_n_3 & ~(sub_666_2_n_2 & n_36));
 assign sub_666_2_n_3 = ~(n_30 & ~n_36);
 assign sub_666_2_n_2 = ~n_30;
 assign sub_666_2_n_1 = ~n_34;
 assign sub_666_2_n_0 = ~n_41;
 assign in2_85_3_ = ~(sub_687_2_n_7 ^ in2_83_2_);
 assign sub_687_2_n_7 = ((sub_687_2_n_5 & sub_687_2_n_0) | ((sub_687_2_n_0 & in2_83_1_) | (in2_83_1_
    & sub_687_2_n_5)));
 assign in2_85_2_ = (sub_687_2_n_0 ^ (in2_83_1_ ^ sub_687_2_n_5));
 assign sub_687_2_n_5 = ((sub_687_2_n_3 & in2_83_0_) | ((in2_83_0_ & sub_687_2_n_1) | (sub_687_2_n_1
    & sub_687_2_n_3)));
 assign in2_85_1_ = (in2_83_0_ ^ (sub_687_2_n_1 ^ sub_687_2_n_3));
 assign in2_85_0_ = ~(sub_687_2_n_3 & ~(sub_687_2_n_2 & n_39));
 assign sub_687_2_n_3 = ~(n_30 & ~n_39);
 assign sub_687_2_n_2 = ~n_30;
 assign sub_687_2_n_1 = ~n_34;
 assign sub_687_2_n_0 = ~n_41;
 assign in2_88_3_ = ~(sub_708_2_n_7 ^ in2_86_2_);
 assign sub_708_2_n_7 = ((sub_708_2_n_5 & sub_708_2_n_0) | ((sub_708_2_n_0 & in2_86_1_) | (in2_86_1_
    & sub_708_2_n_5)));
 assign in2_88_2_ = (sub_708_2_n_0 ^ (in2_86_1_ ^ sub_708_2_n_5));
 assign sub_708_2_n_5 = ((sub_708_2_n_3 & in2_86_0_) | ((in2_86_0_ & sub_708_2_n_1) | (sub_708_2_n_1
    & sub_708_2_n_3)));
 assign in2_88_1_ = (in2_86_0_ ^ (sub_708_2_n_1 ^ sub_708_2_n_3));
 assign in2_88_0_ = ~(sub_708_2_n_3 & ~(sub_708_2_n_2 & n_38));
 assign sub_708_2_n_3 = ~(n_30 & ~n_38);
 assign sub_708_2_n_2 = ~n_30;
 assign sub_708_2_n_1 = ~n_34;
 assign sub_708_2_n_0 = ~n_41;
 assign in2_91_3_ = ~(sub_727_2_n_7 ^ in2_89_2_);
 assign sub_727_2_n_7 = ~((sub_727_2_n_6 | sub_727_2_n_4) & (n_41 | sub_727_2_n_2));
 assign sub_727_2_n_6 = ~((n_28 & sub_727_2_n_3) | (sub_727_2_n_1 & in2_89_0_));
 assign sub_727_2_n_5 = ~({in1[0]} & ~{in2[0]});
 assign sub_727_2_n_4 = ~(in2_89_1_ | ~n_41);
 assign sub_727_2_n_3 = (in2_89_0_ | sub_727_2_n_1);
 assign sub_727_2_n_2 = ~in2_89_1_;
 assign sub_727_2_n_1 = ~n_34;
endmodule

